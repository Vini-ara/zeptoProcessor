library verilog;
use verilog.vl_types.all;
entity Zepto_vlg_vec_tst is
end Zepto_vlg_vec_tst;
