library verilog;
use verilog.vl_types.all;
entity pcTest_vlg_vec_tst is
end pcTest_vlg_vec_tst;
